//0316055_0316313
//Subject:     CO project 3 - Simple Single CPU
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:
//----------------------------------------------
//Date:
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Branch_MUX(
    input branchType_i,
    input zero_i,
    input result_31_i,
    output reg branch_result_o
    );

    

endmodule
